parameter [7:0]  FSIZE = 3;
parameter [7:0]  COF_S = 0;
parameter [7:0]  BPP_S = 1;
