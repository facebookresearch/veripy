parameter   DSS_R1W1   = 0;
parameter   DSS_BE     = 1;
parameter   SYNC_STAGE = 2;

