parameter  DS_X_PP =   2;
parameter  DS_Y_PP =   2;
parameter  PIX_CW  =   11;
parameter  PL      =   10;
parameter  BLOCK   =   3;
parameter  DSXW    =   12;
parameter  NO_RAM  =   BLOCK-1;
parameter  ADDR_W  =   clog2((CAMSIZEX/2)-1);
parameter  PLY     =   5;
parameter  PE      =   5;
parameter  DSY_PP  =   4;
