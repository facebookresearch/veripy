//&module;
module test_verilog_basic1 (
  input  logic        b,
  input  logic        c
); 
//&regs;
//&wires;

wire a = b & c;
endmodule


